netcdf AQUA_MODIS.20020704.L3m.DAY.NSST.sst.4km {
dimensions:
	lat = 4320 ;
	lon = 8640 ;
	rgb = 3 ;
	eightbitcolor = 256 ;
variables:
	short sst(lat, lon) ;
		sst:long_name = "Sea Surface Temperature" ;
		sst:scale_factor = 0.005f ;
		sst:add_offset = 0.f ;
		sst:units = "degree_C" ;
		sst:standard_name = "sea_surface_temperature" ;
		sst:_FillValue = -32767s ;
		sst:valid_min = -1000s ;
		sst:valid_max = 10000s ;
		sst:display_scale = "linear" ;
		sst:display_min = -2.f ;
		sst:display_max = 45.f ;
	ubyte qual_sst(lat, lon) ;
		qual_sst:long_name = "Quality Levels, Sea Surface Temperature" ;
		qual_sst:_FillValue = 255UB ;
		qual_sst:valid_min = 0UB ;
		qual_sst:valid_max = 5UB ;
	float lat(lat) ;
		lat:long_name = "Latitude" ;
		lat:units = "degrees_north" ;
		lat:standard_name = "latitude" ;
		lat:_FillValue = -999.f ;
		lat:valid_min = -90.f ;
		lat:valid_max = 90.f ;
	float lon(lon) ;
		lon:long_name = "Longitude" ;
		lon:units = "degrees_east" ;
		lon:standard_name = "longitude" ;
		lon:_FillValue = -999.f ;
		lon:valid_min = -180.f ;
		lon:valid_max = 180.f ;
	ubyte palette(rgb, eightbitcolor) ;

// global attributes:
		:product_name = "AQUA_MODIS.20020704.L3m.DAY.NSST.sst.4km.nc" ;
		:instrument = "MODIS" ;
		:title = "MODISA Level-3 Standard Mapped Image" ;
		:project = "Ocean Biology Processing Group (NASA/GSFC/OBPG)" ;
		:platform = "Aqua" ;
		:temporal_range = "15-hour" ;
		:processing_version = "R2019.0" ;
		:date_created = "2020-03-19T16:40:13.000Z" ;
		:history = "l3mapgen par=AQUA_MODIS.20020704.L3m.DAY.NSST.sst.4km.nc.param " ;
		:l2_flag_names = "LAND,~HISOLZEN" ;
		:time_coverage_start = "2002-07-04T00:00:10.000Z" ;
		:time_coverage_end = "2002-07-04T14:54:59.000Z" ;
		:start_orbit_number = 885 ;
		:end_orbit_number = 894 ;
		:map_projection = "Equidistant Cylindrical" ;
		:latitude_units = "degrees_north" ;
		:longitude_units = "degrees_east" ;
		:northernmost_latitude = 90.f ;
		:southernmost_latitude = -90.f ;
		:westernmost_longitude = -180.f ;
		:easternmost_longitude = 180.f ;
		:geospatial_lat_max = 90.f ;
		:geospatial_lat_min = -90.f ;
		:geospatial_lon_max = 180.f ;
		:geospatial_lon_min = -180.f ;
		:latitude_step = 0.04166667f ;
		:longitude_step = 0.04166667f ;
		:sw_point_latitude = -89.97916f ;
		:sw_point_longitude = -179.9792f ;
		:spatialResolution = "4.64 km" ;
		:geospatial_lon_resolution = 0.04166667f ;
		:geospatial_lat_resolution = 0.04166667f ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_units = "degrees_east" ;
		:number_of_lines = 4320 ;
		:number_of_columns = 8640 ;
		:measure = "Mean" ;
		:suggested_image_scaling_minimum = -2.f ;
		:suggested_image_scaling_maximum = 45.f ;
		:suggested_image_scaling_type = "LINEAR" ;
		:suggested_image_scaling_applied = "No" ;
		:_lastModified = "2020-03-19T16:40:13.000Z" ;
		:Conventions = "CF-1.6 ACDD-1.3" ;
		:institution = "NASA Goddard Space Flight Center, Ocean Ecology Laboratory, Ocean Biology Processing Group" ;
		:standard_name_vocabulary = "CF Standard Name Table v36" ;
		:naming_authority = "gov.nasa.gsfc.sci.oceandata" ;
		:id = "AQUA_MODIS.20020704.L3b.DAY.NSST.nc/L3/AQUA_MODIS.20020704.L3b.DAY.NSST.nc" ;
		:license = "https://science.nasa.gov/earth-science/earth-science-data/data-information-policy/" ;
		:creator_name = "NASA/GSFC/OBPG" ;
		:publisher_name = "NASA/GSFC/OBPG" ;
		:creator_email = "data@oceancolor.gsfc.nasa.gov" ;
		:publisher_email = "data@oceancolor.gsfc.nasa.gov" ;
		:creator_url = "https://oceandata.sci.gsfc.nasa.gov" ;
		:publisher_url = "https://oceandata.sci.gsfc.nasa.gov" ;
		:processing_level = "L3 Mapped" ;
		:cdm_data_type = "grid" ;
		:data_bins = 3225949LL ;
		:data_minimum = -1.54f ;
		:data_maximum = 32.335f ;
data:

group: processing_control {

  // group attributes:
  		:software_name = "l3mapgen" ;
  		:software_version = "2.3.0-b2c954b" ;
  		:source = "AQUA_MODIS.20020704.L3b.DAY.NSST.nc" ;
  		:l2_flag_names = "LAND,~HISOLZEN" ;

  group: input_parameters {

    // group attributes:
    		:par = "AQUA_MODIS.20020704.L3m.DAY.NSST.sst.4km.nc.param" ;
    		:suite = "NSST" ;
    		:ifile = "AQUA_MODIS.20020704.L3b.DAY.NSST.nc" ;
    		:ofile = "AQUA_MODIS.20020704.L3m.DAY.NSST.sst.4km.nc" ;
    		:oformat = "2" ;
    		:ofile_product_tag = "PRODUCT" ;
    		:ofile2 = "" ;
    		:oformat2 = "png" ;
    		:deflate = "4" ;
    		:product = "sst" ;
    		:resolution = "4km" ;
    		:width = "" ;
    		:projection = "smi" ;
    		:central_meridian = "-999" ;
    		:lat_ts = "" ;
    		:lat_0 = "" ;
    		:lat_1 = "" ;
    		:lat_2 = "" ;
    		:azimuth = "" ;
    		:north = "90.000" ;
    		:south = "-90.000" ;
    		:east = "180.000" ;
    		:west = "-180.000" ;
    		:trimNSEW = "yes" ;
    		:interp = "area" ;
    		:apply_pal = "1" ;
    		:palfile = "" ;
    		:use_transparency = "no" ;
    		:datamin = "" ;
    		:datamax = "" ;
    		:scale_type = "" ;
    		:quiet = "false" ;
    		:pversion = "R2019.0" ;
    		:use_quality = "yes" ;
    		:quality_product = "" ;
    		:use_rgb = "no" ;
    		:product_rgb = "rhos_645,rhos_555,rhos_469" ;
    		:fudge = "1.0" ;
    		:threshold = "0" ;
    		:num_cache = "500" ;
    		:mask_land = "no" ;
    		:land = "$OCDATAROOT/common/landmask_GMT15ARC.nc" ;
    		:full_latlon = "yes" ;
    } // group input_parameters
  } // group processing_control
}
